module FM (
    input wire clk,
    input wire rst_n,
    input wire signed [7:0] d_in,
    input wire [31:0] phi_inc,
    output reg signed [15:0] d_out
);

    wire signed [31:0] port;
    // --- NCO: 单实例同时输出 sin / cos ---
    wire signed [7:0] _nco_sin_u, _nco_cos_u;
    wire signed [15:0] demod_;

    wire signed [7:0] nco_sin, nco_cos;
    assign nco_sin = $signed(_nco_sin_u - 8'd128);
    assign nco_cos = $signed(_nco_cos_u - 8'd128);

    wire signed [15:0] mix_I, mix_Q;

    _NCO #(
    .BASE_PHASE(0)
    ) ncoSin (
        .clk(clk),
        .reset_n(rst_n),
        .phi_inc_i(phi_inc), 
        .nco_out(_nco_sin_u), 
        .out_valid()
    );

    _NCO #(
        .BASE_PHASE(32'h4000_0000) // * 180deg flipped
    ) ncoCos (
        .clk(clk),
        .reset_n(rst_n),
        .phi_inc_i(phi_inc), 
        .nco_out(_nco_cos_u),
        .out_valid()
    );

    // --- Mixing ---
     mixer u_mixer (
        .clk(clk),
        .rst_n(rst_n),
        .adc_data(d_in),
        .nco_sin(nco_sin),  
        .nco_cos(nco_cos),  
        .I_out(mix_I),
        .Q_out(mix_Q)
    );

    // --- FIR Filtering ---
    wire signed [15:0] I_out, Q_out;
    FIR16 fir_I (.clk(clk), .fir_in(mix_I), .fir_out(I_out));
    FIR16 fir_Q (.clk(clk), .fir_in(mix_Q), .fir_out(Q_out));
    // 截断为8位用于后续解调
    wire signed [15:0] I_in = I_out;
    wire signed [15:0] Q_in = Q_out;

    // --- Demodulation (I·Q' - Q·I') ---
    reg signed [15:0] I_prev, Q_prev;
        // 差分处理
    wire signed [15:0] dI = I_in - I_prev;
    wire signed [15:0] dQ = Q_in - Q_prev;
    // demod = I·dQ - Q·dI
    wire signed [31:0] mult1 = I_in * dQ;
    wire signed [31:0] mult2 = Q_in * dI;
    wire signed [31:0] delta_phi = mult1 - mult2;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            I_prev <= 0;
            Q_prev <= 0;
            d_out <= 0;
        end else begin
            I_prev <= I_in;
            Q_prev <= Q_in;
            d_out <= {port[31],port[16:2]}; // 截断为16位输出
        end
    end



    FIR32 fir_demod (.clk(clk), .fir_in(delta_phi), .fir_out(port));

endmodule
