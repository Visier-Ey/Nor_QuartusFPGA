// 63阶 高通FIR滤波器
// 截止频率=0.01π，输入=16位，输出=16位
module FIR_Highpass (
    input clk,
    input signed [15:0] fir_in,
    output signed [15:0] fir_out
);
    reg signed [15:0] delay_line [0:62];

    // 量化系数
    localparam signed [12:0] coeff0 = (-3);
    localparam signed [12:0] coeff1 = (-3);
    localparam signed [12:0] coeff2 = (-3);
    localparam signed [12:0] coeff3 = (-4);
    localparam signed [12:0] coeff4 = (-4);
    localparam signed [12:0] coeff5 = (-5);
    localparam signed [12:0] coeff6 = (-6);
    localparam signed [12:0] coeff7 = (-7);
    localparam signed [12:0] coeff8 = (-8);
    localparam signed [12:0] coeff9 = (-10);
    localparam signed [12:0] coeff10 = (-11);
    localparam signed [12:0] coeff11 = (-13);
    localparam signed [12:0] coeff12 = (-15);
    localparam signed [12:0] coeff13 = (-17);
    localparam signed [12:0] coeff14 = (-19);
    localparam signed [12:0] coeff15 = (-20);
    localparam signed [12:0] coeff16 = (-22);
    localparam signed [12:0] coeff17 = (-24);
    localparam signed [12:0] coeff18 = (-26);
    localparam signed [12:0] coeff19 = (-28);
    localparam signed [12:0] coeff20 = (-30);
    localparam signed [12:0] coeff21 = (-32);
    localparam signed [12:0] coeff22 = (-34);
    localparam signed [12:0] coeff23 = (-35);
    localparam signed [12:0] coeff24 = (-36);
    localparam signed [12:0] coeff25 = (-38);
    localparam signed [12:0] coeff26 = (-39);
    localparam signed [12:0] coeff27 = (-40);
    localparam signed [12:0] coeff28 = (-40);
    localparam signed [12:0] coeff29 = (-41);
    localparam signed [12:0] coeff30 = (-41);
    localparam signed [12:0] coeff31 = (4095);

    always @(posedge clk) begin
        integer i;
        for (i = 62; i > 0; i = i - 1)
            delay_line[i] <= delay_line[i-1];
        delay_line[0] <= fir_in;
    end

    wire signed [28:0] product0, product1, product2, product3, product4, product5, product6, product7, product8, product9, product10, product11, product12, product13, product14, product15, product16, product17, product18, product19, product20, product21, product22, product23, product24, product25, product26, product27, product28, product29, product30, product31;
    assign product0 = (delay_line[0] + delay_line[62]) * coeff0;
    assign product1 = (delay_line[1] + delay_line[61]) * coeff1;
    assign product2 = (delay_line[2] + delay_line[60]) * coeff2;
    assign product3 = (delay_line[3] + delay_line[59]) * coeff3;
    assign product4 = (delay_line[4] + delay_line[58]) * coeff4;
    assign product5 = (delay_line[5] + delay_line[57]) * coeff5;
    assign product6 = (delay_line[6] + delay_line[56]) * coeff6;
    assign product7 = (delay_line[7] + delay_line[55]) * coeff7;
    assign product8 = (delay_line[8] + delay_line[54]) * coeff8;
    assign product9 = (delay_line[9] + delay_line[53]) * coeff9;
    assign product10 = (delay_line[10] + delay_line[52]) * coeff10;
    assign product11 = (delay_line[11] + delay_line[51]) * coeff11;
    assign product12 = (delay_line[12] + delay_line[50]) * coeff12;
    assign product13 = (delay_line[13] + delay_line[49]) * coeff13;
    assign product14 = (delay_line[14] + delay_line[48]) * coeff14;
    assign product15 = (delay_line[15] + delay_line[47]) * coeff15;
    assign product16 = (delay_line[16] + delay_line[46]) * coeff16;
    assign product17 = (delay_line[17] + delay_line[45]) * coeff17;
    assign product18 = (delay_line[18] + delay_line[44]) * coeff18;
    assign product19 = (delay_line[19] + delay_line[43]) * coeff19;
    assign product20 = (delay_line[20] + delay_line[42]) * coeff20;
    assign product21 = (delay_line[21] + delay_line[41]) * coeff21;
    assign product22 = (delay_line[22] + delay_line[40]) * coeff22;
    assign product23 = (delay_line[23] + delay_line[39]) * coeff23;
    assign product24 = (delay_line[24] + delay_line[38]) * coeff24;
    assign product25 = (delay_line[25] + delay_line[37]) * coeff25;
    assign product26 = (delay_line[26] + delay_line[36]) * coeff26;
    assign product27 = (delay_line[27] + delay_line[35]) * coeff27;
    assign product28 = (delay_line[28] + delay_line[34]) * coeff28;
    assign product29 = (delay_line[29] + delay_line[33]) * coeff29;
    assign product30 = (delay_line[30] + delay_line[32]) * coeff30;
    assign product31 = delay_line[31] * coeff31;

    wire signed [34:0] sum = product0 + product1 + product2 + product3 + product4 + product5 + product6 + product7 + product8 + product9 + product10 + product11 + product12 + product13 + product14 + product15 + product16 + product17 + product18 + product19 + product20 + product21 + product22 + product23 + product24 + product25 + product26 + product27 + product28 + product29 + product30 + product31;
    assign fir_out = sum[34:19];
endmodule