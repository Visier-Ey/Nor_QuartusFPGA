`timescale 1us/1us

module touch_led_tb();


touch_key u_touch_key(){
    
}

endmodule